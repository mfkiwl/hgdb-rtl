module mod1;
endmodule;

module top;
mod1 inst0();
mod1 inst1();
mod1 inst12();
endmodule
